`timescale 1ns/10ps

module alu_test;
	reg		[31:0]	A, B;
	reg		[3:0] 	ctrl;
	wire 			cout, over, zero;
	wire	[31:0]	res;
	 
	alu alu0(A, B, ctrl, cout, over, zero, res);
	
	initial $monitor ("A: %d B: %d      cout: %b over: %b zero: %b res: %d", 
						$signed(A), $signed(B), cout, over, zero, $signed(res));

	integer i;

// insert data
	initial 
		begin
// Test add
			$display("--------------------------------------------");
			$display("Test Add");
			ctrl = 4'b0010;
// 0 + 0
			A = 0;
			B = 0;
			#10
// 0 + 100
			A = 0;
			B = 100;
			#10
// 100 + 0
			A = 100;
			B = 0;
			#10
// 100 + 100
			A = 100;
			B = 100;
			#10
// 2147483647 + 0
			A = 2147483647;
			B = 0;
			#10
// 1 + 2147483647 OVERFLOW
			A = 1;
			B = 2147483647;
			#10
// -1 + 1 CARRY OUT
			A = -1;
			B = 1;
			#20



// Test sub
			$display("--------------------------------------------");
			$display("Test Sub");
			ctrl = 4'b0110;
// 0 - 0
			A = 0;
			B = 0;
			#10
// -1 - -1
			A = -1;
			B = -1;
			#10
// 0 - 100
			A = 0;
			B = 100;
			#10
// 100 - 0
			A = 100;
			B = 0;
			#10
// 100 - 100
			A = 100;
			B = 100;
			#10
// 100 - 99
			A = 100;
			B = 99;
			#10	
// 2147483647 - -1 OVERFLOW
			A = 2147483647;
			B = -1;
			#10	
// -2147483648 - 1 UNDERFLOW
			A = -2147483648;
			B = 1;
			#10	
// 1 - 2	UNSIGNED CARRYOUT 0
			A = 1;
			B = 2;
			#20



// Test and 
			$display("--------------------------------------------");
			$display("Test And");
			ctrl = 4'b0000;
// 0 and 0
			A = 0;
			B = 0;
			#10
// -1 and 0
			A = -1;
			B = 0;
			#10
// 0 and -1
			A = 0;
			B = -1;
			#10
// -1 and -1
			A = -1;
			B = -1;
			#10
// 99 and 100 = 96
			A = 99;
			B = 100;
			#20



// Test or 
			$display("--------------------------------------------");
			$display("Test Or");
			ctrl = 4'b0001;
// 0 and 0
			A = 0;
			B = 0;
			#10
// -1 and 0
			A = -1;
			B = 0;
			#10
// 0 and -1
			A = 0;
			B = -1;
			#10
// -1 and -1
			A = -1;
			B = -1;
			#10
// 99 and 100 = 103
			A = 99;
			B = 100;
			#20



// Test xor 
			$display("--------------------------------------------");
			$display("Test Xor");
			ctrl = 4'b0011;
// 0 and 0
			A = 0;
			B = 0;
			#10
// -1 and 0
			A = -1;
			B = 0;
			#10
// 0 and -1
			A = 0;
			B = -1;
			#10
// -1 and -1
			A = -1;
			B = -1;
			#10
// 99 and 100 = 7
			A = 99;
			B = 100;
			#20

			

// Test SLT 
			$display("--------------------------------------------");
			$display("Test slt");
			ctrl = 4'b0111;
// 0 < 100
			A = 0;
			B = 100;
			#10
// -1 < 100
			A = -1;
			B = 100;
			#10
// -1 < 0
			A = -1;
			B = 0;
			#10
// 0 < 0
			A = 0;
			B = 0;
			#10
// -1 < -1
			A = -1;
			B = -1;
			#10
// 0 < -1
			A = 0;
			B = -1;
			#10
// -1 < -2147483648
			A = -1;
			B = -2147483648;
			#10
// -3 < -2147483648
			A = -3;
			B = -2147483648;
			#10
// -2147483648 < -2147483648
			A = -2147483648;
			B = -2147483648;
			#10
// -2147483647 < -2147483648
			A = -2147483647;
			B = -2147483648;
			#10
// -2147483648 < -2147483647
			A = -2147483648;
			B = -2147483647;
			#10
// 1 < 2147483647
			A = 1;
			B = 2147483647;
			#10
// 2147483647 < 2147483647
			A = 2147483647;
			B = 2147483647;
			#10
// 2147483646 < 2147483647
			A = 2147483646;
			B = 2147483647;
// -2147483648 < 2147483647
			A = -2147483648;
			B = 2147483647;
			#20



// Test SLTU 
			$display("--------------------------------------------");
			$display("Test Sltu");
			ctrl = 4'b0101;
		
// 0 < 100
			A = 0;
			B = 100;
			#10
// 0 < 0
			A = 0;
			B = 0;
			#10
// -1 < 0
			A = -1;
			B = 0;
			#10
// 0 < -1
			A = 0;
			B = -1;
			#10
// -2 < -1
			A = -2;
			B = -1;
			#10
// -1 < -2
			A = -1;
			B = -2;
			#10
// 999 < 1000
			A = 999;
			B = 1000;
			#10
// 1000 < 999
			A = 1000;
			B = 999;
			#10
// -100 < -99
			A = -100;
			B = -99;
			#10
// -999 < -999
			A = -999;
			B = -999;
			#10
// -99 < -100
			A = -99;
			B = -100;
			#20

// Test Left Shift
			$display("--------------------------------------------");
			$display("Test Left Shift");
			ctrl = 4'b1000;

			A = 32'b01010101010101010101010101010101; 
			for (i = 0; i < 32; i = i + 1) begin
				B = i;
				#1;
			end
			#10

			$display("\n\n");
			A = 32'b10101010101010101010101010101010; 
			for (i = 0; i < 32; i = i + 1) begin
				B = i;
				#1;
			end

// Test Right Shift
			$display("--------------------------------------------");
			$display("Test Right Shift");
			ctrl = 4'b1001;

			A = 32'b01010101010101010101010101010101; 
			for (i = 0; i < 32; i = i + 1) begin
				B = i;
				#1;
			end
			#10

			$display("\n\n");
			A = 32'b10101010101010101010101010101010; 
			for (i = 0; i < 32; i = i + 1) begin
				B = i;
				#1;
			end

// Test random
			$display("--------------------------------------------");
			$display("Test Random");
			ctrl = 4'b0010;
			A = 32'h00afb000;
			B = -32'h000f0000;
			#10

			ctrl = 4'b0000;
			A = 32'hff00f00f;
			B = 32'h1f00100f;
			#10

            #20 $finish;
			
	end 
endmodule
